* ---------- MODEL 1 ----------
.MODEL MODEL1 NPN (IS=10e-15 BF=200 XTI=3E00 VAR=1.00E2 IKF=46.7E-03
+EG=1.110E00 VAF=150 ISE=114.286E-15 NE=1.48E00 XTB=0
+BR=0.1 ISC=10.005e-15 NC=2 IKR=10e-3 RC=10 
+MJC=.333 VJC=.75 FC=5.00e-01 CJE=1.02e-12 MJE=.336 VJE=.75
+TR=10e-9 TF=277.01e-12 ITF=1.75 XTF=309.38 VTF=16.37)

* ---------- MODEL 2 ----------
.MODEL MODEL2 NPN (IS=10e-15 BF=150 XTI=3E00 VAR=1.00E2 IKF=46.7E-03
+EG=1.110E00 VAF=120 ISE=114.286E-15 NE=1.48E00 XTB=0
+BR=0.1 ISC=10.005e-15 NC=2 IKR=10e-3 RC=10 
+MJC=.333 VJC=.75 FC=5.00e-01 CJE=1.02e-12 MJE=.336 VJE=.75
+TR=10e-9 TF=277.01e-12 ITF=1.75 XTF=309.38 VTF=16.37)

* ---------- MODEL 3 ----------
.MODEL MODEL3 NPN (IS=10e-15 BF=100 XTI=3E00 VAR=1.00E2 IKF=46.7E-03
+EG=1.110E00 VAF=100 ISE=114.286E-15 NE=1.48E00 XTB=0
+BR=0.1 ISC=10.005e-15 NC=2 IKR=10e-3 RC=10 
+MJC=.333 VJC=.75 FC=5.00e-01 CJE=1.02e-12 MJE=.336 VJE=.75
+TR=10e-9 TF=277.01e-12 ITF=1.75 XTF=309.38 VTF=16.37)

* ---------- MODEL 4 ----------
.MODEL MODEL4 NPN (IS=10e-15 BF=80 XTI=3E00 VAR=1.00E2 IKF=46.7E-03
+EG=1.110E00 VAF=80 ISE=114.286E-15 NE=1.48E00 XTB=0
+BR=0.1 ISC=10.005e-15 NC=2 IKR=10e-3 RC=10 
+MJC=.333 VJC=.75 FC=5.00e-01 CJE=1.02e-12 MJE=.336 VJE=.75
+TR=10e-9 TF=277.01e-12 ITF=1.75 XTF=309.38 VTF=16.37)

* ---------- MODEL 5 ----------
.MODEL MODEL5 NPN (IS=10e-15 BF=50 XTI=3E00 VAR=1.00E2 IKF=46.7E-03
+EG=1.110E00 VAF=50 ISE=114.286E-15 NE=1.48E00 XTB=0
+BR=0.1 ISC=10.005e-15 NC=2 IKR=10e-3 RC=10 
+MJC=.333 VJC=.75 FC=5.00e-01 CJE=1.02e-12 MJE=.336 VJE=.75
+TR=10e-9 TF=277.01e-12 ITF=1.75 XTF=309.38 VTF=16.37)
