* MODEL 1
.model MODEL1 NPN (BF=200 VAF=1000 IS=1e-15)

* MODEL 2
.model MODEL2 NPN (BF=150 VAF=1000 IS=1e-15)

* MODEL 3
.model MODEL3 NPN (BF=120 VAF=1000 IS=1e-15)

*MODEL 4
.model MODEL4 NPN (BF=100 VAF=1000 IS=1e-15)

*MODEL 5
.model MODEL5 NPN (BF=80 VAF=1000 IS=1e-15)