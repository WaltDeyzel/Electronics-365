*------------------------------------------------------------------------------------------------------------------------- * SPICE model for amplifier with compensation
* -------------------------------------------
* Surname: Your surname
* First name: Your first name
* Student number: Your student number
* -------------------------------------------

* op amp model
.subckt opamp   non    inv     out
Ri      non    inv     1e14
Eout    out    0       non    inv    1e7
.ends

* Define amplifier circuit with compensation as a subcircuit
.subckt comps pa na pb nb vcc vee vo1 vo2 vx1 vx2

* -------- Start of student code --------

*Op amps for amplifier
XOPAMPA  pa   na   vo1   opamp
XOPAMPB  pb   nb   vo2   opamp

* Original circuit with random values
R1      0     na     20k
R2      na    vo1    80k
R3      vx3   nb     15k
R4      nb    vo2    45k

* Dummy components in the place of compensation
Rd1  pa  0    16k
Rd2  pb   pb  11.25k
Rd3  vx3  0    11k

* --------- End of student code ---------
.ends
*-------------------------------------------------------------------------------------------------------------------------
