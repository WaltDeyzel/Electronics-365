*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Inc.
* Models developed and under copyright by:
* National Semiconductor, Inc.

*/////////////////////////////////////////////////////////////////////
* Legal Notice: This material is intended for free software support.
* The file may be copied, and distributed; however, reselling the
*  material is illegal

*////////////////////////////////////////////////////////////////////
* For ordering or technical information on these models, contact:
* National Semiconductor's Customer Response Center
*                 7:00 A.M.--7:00 P.M.  U.S. Central Time
*                                (800) 272-9959
* For Applications support, contact the Internet address:
*  amps-apps@galaxy.nsc.com

*//////////////////////////////////////////////////////////
*LM741 OPERATIONAL AMPLIFIER MACRO-MODEL
*//////////////////////////////////////////////////////////
*
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   positive power supply
*                   |   |   |   negative power supply
*                   |   |   |   |   output
*                   |   |   |   |   |
*                   |   |   |   |   |
.SUBCKT LM741/NS    1   2  99  50  28
*
*Features:
*Improved performance over industry standards
*Plug-in replacement for LM709,LM201,MC1439,748
*Input and output overload protection
*
****************INPUT STAGE**************
*
IOS 2 1 20N
*^Input offset current
R1 1 3 250K
R2 3 2 250K
I1 4 50 100U
R3 5 99 517
R4 6 99 517
Q1 5 2 4 QX
Q2 6 7 4 QX
*Fp2=2.55 MHz
C4 5 6 60.3614P
*
***********COMMON MODE EFFECT***********
*
I2 99 50 1.6MA
*^Quiescent supply current
EOS 7 1 POLY(1) 16 49 1E-3 1
*Input offset voltage.^
R8 99 49 40K
R9 49 50 40K
*
*********OUTPUT VOLTAGE LIMITING********
V2 99 8 1.63
D1 9 8 DX
D2 10 9 DX
V3 10 50 1.63
*
**************SECOND STAGE**************
*
EH 99 98 99 49 1
G1 98 9 5 6 2.1E-3
*Fp1=5 Hz
R5 98 9 95.493MEG
C3 98 9 333.33P
*
***************POLE STAGE***************
*
*Fp=30 MHz
G3 98 15 9 49 1E-6
R12 98 15 1MEG
C5 98 15 5.3052E-15
*
*********COMMON-MODE ZERO STAGE*********
*
*Fpcm=300 Hz
G4 98 16 3 49 3.1623E-8
L2 98 17 530.5M
R13 17 16 1K
*
**************OUTPUT STAGE**************
*
F6 50 99 POLY(1) V6 450U 1
E1 99 23 99 15 1
R16 24 23 25
D5 26 24 DX
V6 26 22 0.65V
R17 23 25 25
D6 25 27 DX
V7 22 27 0.65V
V5 22 21 0.18V
D4 21 15 DX
V4 20 22 0.18V
D3 15 20 DX
L3 22 28 100P
RL3 22 28 100K
*
***************MODELS USED**************
*
.MODEL DX D(IS=1E-15)
.MODEL QX NPN(BF=625)
*
.ENDS
*$
****************************************
*Section A circuit
Vcc     vcc    0    DC    15
Vee     vee    0    DC   -15

XopampA  ni      in  vcc    vee    out    LM741/NS

R1      xxx    in  2k
R2      inv   out  8k
r		ni     0    0
RL      out    0    150k

vi      111    0    0    ac    1    0
Rs      111    xxx  50

.control
   * Do AC sweep when AvCL approxeq 1E6
  AC    DEC   101   1   10E6
   * Result available in ac1.
   * Now change resistance of R2 to 100000 kOhm; AvCL = 1E5
  *alter @r2[r]=100000k
   * Do the AC sweep for AvCL = 1E5
  *AC    DEC   101   1   10E6
   * Result available in ac2.
   * Now change resistance of R2 to 10000 kOhm; AvCL = 1E4
  *alter @r2[r]=10000k
  *AC    DEC   101   1   10E6
   * Result in ac3. Repeat pattern: R2 changed to 1000 kOhm
  *alter @r2[r]=1000k
  *AC    DEC   101   1   10E6
  *alter @r2[r]=100k
  *AC    DEC   101   1   10E6
  *alter @r2[r]=10k
  *AC    DEC   101   1   10E6
  *alter @r2[r]=1k
  *AC    DEC   101   1   10E6


   * Calculate gain vs frequency in dB fro ac1
  let  run1db = 20*log10(abs(ac1.v(out)))
   * And do for the other runs too
  *let  run2db = 20*log10(abs(ac2.v(out)))
  *let  run3db = 20*log10(abs(ac3.v(out)))
  *let  run4db = 20*log10(abs(ac4.v(out)))
  *let  run5db = 20*log10(abs(ac5.v(out)))
  *let  run6db = 20*log10(abs(ac6.v(out)))
  *let  run7db = 20*log10(abs(ac7.v(out)))

   * Plot all on the same plot
  plot run1db
*run2db run3db run4db run5db run6db run7db
.endc

.end
